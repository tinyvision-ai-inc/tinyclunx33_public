`define FAST_SIM